module TSC (
  input wire clk 
);
endmodule

